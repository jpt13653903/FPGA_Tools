//==============================================================================
// Copyright (C) John-Philip Taylor
// jpt13653903@gmail.com
//
// This file is part of a library
//
// This file is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>
//==============================================================================

// n-bit synchronous up-counter

module Counter #(
  parameter n = 8
)(
  input nReset, 
  input Clk, 

  output reg [n-1:0]Output
);
//------------------------------------------------------------------------------
 
  always @(negedge nReset, negedge Clk) begin
    if(!nReset) Output <= 0;
    else        Output <= Output + 1'b1;
  end
endmodule
//------------------------------------------------------------------------------

