//==============================================================================
// Copyright (C) John-Philip Taylor
// jpt13653903@gmail.com
//
// This file is part of S/PDIF Radio
//
// This file is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>
//==============================================================================

module SD_Data_Bus #(
  parameter Bus_Width = 4 // Either 1 or 4
)(
  input Reset,
  input Clk,    // Controller clock
  input SD_Clk, // The SD-Card clock, generated by the controller.  The real
                // clock (output to the SD-card) is delayed by one Clk cycle.

  input [11:0]Block_Length, // N-1, per data line, excluding CRC and admin
  input       Send,         // Starts a send cycle, 
                            // receiving starts automatically on a start bit

  output reg      Data_Clk,  // Controls the data stream, data is read / written 
  output reg [7:0]Receive_Data, // on every edge
  input      [7:0]Send_Data,

  output reg      Busy,  // High while busy sending / receiving
  output reg [3:0]Error, // Used for both send and receive upon CRC fail

  inout  reg [3:0]SD_Data,
  output          SD_Busy // Sampled on the correct edge
);
//------------------------------------------------------------------------------

assign SD_Busy = ~tSD_Data[0];
//------------------------------------------------------------------------------

// States:
reg   [2:0]State;
localparam Idle         = 3'b000;
localparam Sending      = 3'b001;
localparam SendingCRC   = 3'b011;
localparam Response     = 3'b010; // Get CRC and busy response from card
localparam Done         = 3'b110;

localparam Receiving    = 3'b100;
localparam ReceivingCRC = 3'b101;

integer j;

reg      pSD_Clk;
reg [3:0]tSD_Data;

reg [11:0]Count;
reg [15:0]CRC   [3:0];
reg [15:0]CRC_In[3:0];
reg [ 6:0]Temp;
//------------------------------------------------------------------------------

reg tReset;

always @(posedge Clk) begin
  tReset <= Reset;

  if(tReset) begin
    State   <= Idle;
    pSD_Clk <= 0;

    Data_Clk     <= 0;
    Receive_Data <= 0;
    Busy         <= 0;
    Error        <= 0;
    SD_Data      <= 4'bZZZZ;
    tSD_Data     <= 4'b1111;

    Count     <= 0;
    CRC   [0] <= 0;
    CRC   [1] <= 0;
    CRC   [2] <= 0;
    CRC   [3] <= 0;
    CRC_In[0] <= 0;
    CRC_In[1] <= 0;
    CRC_In[2] <= 0;
    CRC_In[3] <= 0;
    Temp      <= 0;
//------------------------------------------------------------------------------
  
  end else begin
    pSD_Clk <= SD_Clk;
//------------------------------------------------------------------------------

    if(pSD_Clk & ~SD_Clk) begin // Falling edge (host to card)
      if(Bus_Width == 4) tSD_Data <=          SD_Data;
      else               tSD_Data <= {3'b111, SD_Data[0]};

      case(State)
        Idle: begin
          if(Send) begin
            Busy  <= 1'b1;
            Error <= 4'd0;
            State <= Done;
          end
        end
//------------------------------------------------------------------------------

        Sending: begin
        end
//------------------------------------------------------------------------------

        SendingCRC: begin
        end
//------------------------------------------------------------------------------

        Response: begin
        end
//------------------------------------------------------------------------------

        Done: begin
          if(~Send) begin
            Busy  <= 1'b0;
            State <= Idle;
          end
        end
//------------------------------------------------------------------------------

        default:;
      endcase;
//------------------------------------------------------------------------------

    end else if(~pSD_Clk & SD_Clk) begin // Rising edge (card to host)
      case(State)
        Idle: begin
          if(~&tSD_Data) begin
            Count  <= Block_Length;
            CRC[0] <= 16'd0;
            CRC[1] <= 16'd0;
            CRC[2] <= 16'd0;
            CRC[3] <= 16'd0;
            Busy   <=  1'b1;
            Error  <=  4'd0;
            State  <= Receiving;
          end
        end
//------------------------------------------------------------------------------

        Receiving: begin
          if(Bus_Width == 4) begin
            if(Count[0]) begin
              Temp[3:0] <= tSD_Data;
            end else begin
              Data_Clk     <= ~Data_Clk;
              Receive_Data <= {Temp[3:0], tSD_Data};
            end
          end else begin
            if(|Count[2:0]) begin
              Temp <= {Temp[5:0], tSD_Data[0]};
            end else begin
              Data_Clk     <= ~Data_Clk;
              Receive_Data <= {Temp, tSD_Data[0]};
            end
          end

          for(j = 0; j < Bus_Width; j = j + 1) begin
            CRC[j] <= {
              CRC[j][14:12], 
              CRC[j][   11]^ (tSD_Data[j] ^ CRC[j][15]),
              CRC[j][10: 5], 
              CRC[j][    4]^ (tSD_Data[j] ^ CRC[j][15]),
              CRC[j][ 3: 0], (tSD_Data[j] ^ CRC[j][15])
            };
          end

          if(~|Count) begin
            Count[4:0] <= 5'd16;
            State <= ReceivingCRC;
          end else begin
            Count <= Count - 1'b1;
          end
        end
//------------------------------------------------------------------------------

        ReceivingCRC: begin
          for(j = 0; j < Bus_Width; j = j + 1) begin
            CRC_In[j] <= {CRC_In[j][14:0], tSD_Data[j]};
          end

          if(~|Count[4:0]) begin
            Error[0] <= (CRC[0] != CRC_In[0]);
            if(Bus_Width == 4) begin
              Error[1] <= (CRC[1] != CRC_In[1]);
              Error[2] <= (CRC[2] != CRC_In[2]);
              Error[3] <= (CRC[3] != CRC_In[3]);
            end else begin
              Error[1] <= 1'b0;
              Error[2] <= 1'b0;
              Error[3] <= 1'b0;
            end
            Busy  <= 1'b0;
            State <= Idle;

          end else begin
            Count[4:0] <= Count[4:0] - 1'b1;
          end
        end
//------------------------------------------------------------------------------

        default:;
      endcase
    end  
  end
end
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

