`define ALU_Add         4'd0
`define ALU_And         4'd1
`define ALU_Or          4'd2
`define ALU_XOr         4'd3
`define ALU_RotateLeft  4'd4
`define ALU_RotateRight 4'd5
`define ALU_Swap        4'd6
`define ALU_BitSet      4'd7
`define ALU_BitClear    4'd8
`define ALU_BitTest     4'd9

