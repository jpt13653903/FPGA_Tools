--==============================================================================
-- Copyright (C) John-Philip Taylor
-- jpt13653903@gmail.com
--
-- This file is part of a library
--
-- This file is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>
--==============================================================================

-- J Taylor
-- Last modified 2009-11-23
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--------------------------------------------------------------------------------

entity CPU_Adder is
 port(
  A        : in  std_logic_vector(7 downto 0);
  B        : in  std_logic_vector(8 downto 0);
  Carry_In : in  std_logic;
  Y        : out std_logic_vector(7 downto 0);
  Carry    : out std_logic
 );
end entity CPU_Adder;
--------------------------------------------------------------------------------

architecture a1 of CPU_Adder is
 signal tY : std_logic_vector(8 downto 0);
begin
 tY     <= A + B + Carry_In;
 Y      <= tY(7 downto 0);
 Carry  <= tY(8);
end architecture a1;
--------------------------------------------------------------------------------
